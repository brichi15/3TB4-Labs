module test (x,q);


endmodule